// Memory for Multi-cycle Implementation

module Memory(MemData,Address,WriteData,MemRead,MemWrite,Clock);

   // Port Declarations
   output [31:0] MemData;
   input [31:0]  WriteData,Address; 
   input 	 MemRead,MemWrite,Clock;

   reg [7:0] 	 Memory[0:1023];

   initial
     begin
	//ADD Rd,Rs1,Rs2 000000 10001 10010 00001 00000 000100
	{Memory[0],Memory[1],Memory[2],Memory[3]} = 32'b000000_10000_10010_00001_00000_000100;
	//SUB Rd,Rs1,Rs2 000000 10001 10010 00001 00000 000110
	{Memory[4],Memory[5],Memory[6],Memory[7]} = 32'b000000_10001_10010_00001_00000_000110;
	//AND Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001000
	{Memory[8],Memory[9],Memory[10],Memory[11]} = 32'b000000_10001_10010_00001_00000_001000;
	//OR  Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001001
	{Memory[12],Memory[13],Memory[14],Memory[15]} = 32'b000000_10001_10010_00001_00000_001001;
	//XOR Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001010
	{Memory[16],Memory[17],Memory[18],Memory[19]} = 32'b000000_10001_10010_00001_00000_001010;
	//SLL Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001100
	{Memory[20],Memory[21],Memory[22],Memory[23]} = 32'b000000_10001_10010_00001_00000_001100;
	//SRL Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001110
	{Memory[24],Memory[25],Memory[26],Memory[27]} = 32'b000000_10001_10010_00001_00000_001110;
	//SRA Rd,Rs1,Rs2 000000 10001 10010 00001 00000 001111
	{Memory[28],Memory[29],Memory[30],Memory[31]} = 32'b000000_10001_10010_00001_00000_001111;

	//I
	//ADDI Rd,Rs1,Imm 010100 10001 00001 0000000011001100 204
	{Memory[32],Memory[33],Memory[34],Memory[35]} = 32'b010100_10001_00001_0000000011001100;
	//SUBI Rd,Rs1,Imm 010110 10001 00001 0000000011001100
	{Memory[36],Memory[37],Memory[38],Memory[39]} = 32'b010110_10001_00001_0000000011001100;
	//ANDI Rd,Rs1,Imm 011000 10001 00001 0000000011001100
	{Memory[40],Memory[41],Memory[42],Memory[43]} = 32'b011000_10001_00001_0000000011001100;
	//ORI  Rd,Rs1,Imm 011001 10001 00001 0000000011001100
	{Memory[44],Memory[45],Memory[46],Memory[47]} = 32'b011001_10001_00001_0000000011001100;
	//XORI Rd,Rs1,Imm 011010 10001 00001 0000000011001100
	{Memory[48],Memory[49],Memory[50],Memory[51]} = 32'b011010_10001_00001_0000000011001100;
	//SLLI Rd,Rs1,Imm 011100 10001 00001 0000000011001100
	{Memory[52],Memory[53],Memory[54],Memory[55]} = 32'b011100_10001_00001_0000000011001100;
	//SRLI Rd,Rs1,Imm 011110 10001 00001 0000000011001100
	{Memory[56],Memory[57],Memory[58],Memory[59]} = 32'b011110_10001_00001_0000000011001100;
	//SRAI Rd,Rs1,Imm 011111 10001 00001 0000000011001100
	{Memory[60],Memory[61],Memory[62],Memory[63]} = 32'b011111_10001_00001_0000000011001100;
	//LHI  Rd,Rs1,Imm 011011 10001 00001 0000000011001100
	{Memory[64],Memory[65],Memory[66],Memory[67]} = 32'b011011_10001_00001_0000000011001100;

	//NOP Rd,Rs1,Rs2 000000 00000 00000 00000 00000 000000
	{Memory[68],Memory[69],Memory[70],Memory[71]} = 32'b000000_00000_00000_00000_00000_000000;
	//SEQ Rd,Rs1,Rs2 000000 10001 10010 00001 00000 010000
	{Memory[72],Memory[73],Memory[74],Memory[75]} = 32'b000000_10001_10010_00001_00000_010000;
	//SNE Rd,Rs1,Rs2 000000 10001 10010 00001 00000 010010
	{Memory[76],Memory[77],Memory[78],Memory[79]} = 32'b000000_10001_10010_00001_00000_010010;
	//SLT Rd,Rs1,Rs2 000000 10001 10010 00001 00000 010100
	{Memory[80],Memory[81],Memory[82],Memory[83]} = 32'b000000_10001_10010_00001_00000_010100;
	//SLE Rd,Rs1,Rs2 000000 10001 10010 00001 00000 010110
	{Memory[84],Memory[85],Memory[86],Memory[87]} = 32'b000000_10001_10010_00001_00000_010110;
	//SGT Rd,Rs1,Rs2 000000 10001 10010 00001 00000 011000
	{Memory[88],Memory[89],Memory[90],Memory[91]} = 32'b000000_10001_10010_00001_00000_011000;
	//SGE Rd,Rs1,Rs2 000000 10001 10010 00001 00000 011010
	{Memory[92],Memory[93],Memory[94],Memory[95]} = 32'b000000_10001_10010_00001_00000_011010;

	//I
	//SEQI  Rd,Rs1,Imm 100000 10001 00001 0000000011001100
	{Memory[96],Memory[97],Memory[98],Memory[99]} = 32'b100000_10001_00001_0000000011001100;
	//SNEI  Rd,Rs1,Imm 100010 10001 00001 0000000011001100
	{Memory[100],Memory[101],Memory[102],Memory[103]} = 32'b100010_10001_00001_0000000011001100;
	//SLTI  Rd,Rs1,Imm 100100 10001 00001 0000000011001100
	{Memory[104],Memory[105],Memory[106],Memory[107]} = 32'b100100_10001_00001_0000000011001100;
	//SLEI  Rd,Rs1,Imm 100110 10001 00001 0000000011001100
	{Memory[108],Memory[109],Memory[110],Memory[111]} = 32'b100110_10001_00001_0000000011001100;
	//SGTI  Rd,Rs1,Imm 101000 10001 00001 0000000011001100
	{Memory[112],Memory[113],Memory[114],Memory[115]} = 32'b101000_10001_00001_0000000011001100;
	//SGEI  Rd,Rs1,Imm 101010 10001 00001 0000000011001100
	{Memory[116],Memory[117],Memory[118],Memory[119]} = 32'b101010_10001_00001_0000000011001100;
	
     end // initial begin

   // Read from memory
   assign MemData = MemRead ? {Memory[Address],Memory[Address+1],Memory[Address+2],Memory[Address+3]} :0;

   //Write to memory
   always @ (posedge Clock) 
     begin
	if (MemWrite) 
	  begin
	     Memory[Address] <= WriteData; 
	  end
     end
endmodule // Memory
